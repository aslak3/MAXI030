`define TIMER_INT_POS   0
`define QUART_INT_POS   1
`define IDE_INT_POS     2
`define ETH_INT_POS     3
`define PS2_INT_POS     4
